module q_sys_pll_status_interconnect_2 (
		input  wire [0:0] pll_locked,        //        pll_locked.pll_locked
		output wire [0:0] pll_powerdown,     //     pll_powerdown.pll_powerdown
		output wire [0:0] mcgb_rst,          //          mcgb_rst.mcgb_rst
		output wire [0:0] pll_locked_output, // pll_locked_output.pll_locked
		output wire [0:0] pll_locked_a,      //      pll_locked_a.pll_locked
		input  wire [0:0] pll_powerdown_a,   //   pll_powerdown_a.pll_powerdown
		output wire [0:0] pll_locked_b,      //      pll_locked_b.pll_locked
		input  wire [0:0] pll_powerdown_b    //   pll_powerdown_b.pll_powerdown
	);
endmodule

