module q_sys_clock_bridge_1 (
		input  wire  in_clk,  //  in_clk.clk
		output wire  out_clk  // out_clk.clk
	);
endmodule

