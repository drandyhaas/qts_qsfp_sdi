module sdi_xcvr_test_clk_100 (
		input  wire  in_clk,      //       clk_in.clk
		input  wire  reset_n,     // clk_in_reset.reset_n
		output wire  clk_out,     //          clk.clk
		output wire  reset_n_out  //    clk_reset.reset_n
	);
endmodule

