module xcvr_test_system_xcvr_tx_rx_clkout2_converter_0 (
		input  wire  rx_clkout2,        //        rx_clkout2.clk
		output wire  rx_clkout2_a,      //      rx_clkout2_a.export
		output wire  rx_clkout2_b,      //      rx_clkout2_b.export
		input  wire  tx_clkout2,        //        tx_clkout2.clk
		output wire  tx_clkout2_a,      //      tx_clkout2_a.export
		output wire  tx_clkout2_b,      //      tx_clkout2_b.export
		output wire  tx_clkout2_sample  // tx_clkout2_sample.clk
	);
endmodule

