// qsfp_xcvr_test.v

// Generated using ACDS version 23.3 104

`timescale 1 ps / 1 ps
module qsfp_xcvr_test (
		input  wire        clk_100_clk,                                     //                          clk_100.clk
		input  wire        reset_100_reset_n,                               //                        reset_100.reset_n
		input  wire        clk_50_clk,                                      //                           clk_50.clk
		input  wire        reset_50_reset_n,                                //                         reset_50.reset_n
		output wire        mm_bridge_0_s0_waitrequest,                      //                   mm_bridge_0_s0.waitrequest
		output wire [31:0] mm_bridge_0_s0_readdata,                         //                                 .readdata
		output wire        mm_bridge_0_s0_readdatavalid,                    //                                 .readdatavalid
		input  wire [0:0]  mm_bridge_0_s0_burstcount,                       //                                 .burstcount
		input  wire [31:0] mm_bridge_0_s0_writedata,                        //                                 .writedata
		input  wire [14:0] mm_bridge_0_s0_address,                          //                                 .address
		input  wire        mm_bridge_0_s0_write,                            //                                 .write
		input  wire        mm_bridge_0_s0_read,                             //                                 .read
		input  wire [3:0]  mm_bridge_0_s0_byteenable,                       //                                 .byteenable
		input  wire        mm_bridge_0_s0_debugaccess,                      //                                 .debugaccess
		input  wire [0:0]  pll_locked_pll_locked_pll_locked,                //            pll_locked_pll_locked.pll_locked
		input  wire [0:0]  xcvr_native_s10_0_tx_serial_clk0_clk,            // xcvr_native_s10_0_tx_serial_clk0.clk
		input  wire        xcvr_native_s10_0_rx_cdr_refclk0_clk,            // xcvr_native_s10_0_rx_cdr_refclk0.clk
		output wire [0:0]  xcvr_native_s10_0_tx_serial_data_tx_serial_data, // xcvr_native_s10_0_tx_serial_data.tx_serial_data
		input  wire [0:0]  xcvr_native_s10_0_rx_serial_data_rx_serial_data  // xcvr_native_s10_0_rx_serial_data.rx_serial_data
	);

	wire         clk_50_clk_clk;                                                                             // clk_50:clk_out -> [default_pma_settings_conf_0:clock, mm_bridge_0:clk, mm_interconnect_0:clk_50_clk_clk, nativePHY_loopback_cont_0:clk, rst_controller:clk, xcvr_test_system_0:clk_50_clk]
	wire         clk_100_clk_clk;                                                                            // clk_100:clk_out -> [mm_interconnect_0:clk_100_clk_clk, rst_controller_001:clk, xcvr_native_s10_0:reconfig_clk, xcvr_reset_control_s10_0:clock]
	wire   [0:0] xcvr_native_s10_0_rx_clkout_clk;                                                            // xcvr_native_s10_0:rx_clkout -> xcvr_st_converter_0:rx_clkout
	wire   [0:0] xcvr_native_s10_0_rx_clkout2_clk;                                                           // xcvr_native_s10_0:rx_clkout2 -> xcvr_test_system_0:xcvr_tx_rx_clkout2_converter_0_rx_clkout2_clk
	wire         xcvr_st_converter_0_rx_clkout_a_output_clk;                                                 // xcvr_st_converter_0:rx_clkout_a_output -> xcvr_native_s10_0:rx_coreclkin
	wire   [0:0] xcvr_native_s10_0_tx_clkout_clk;                                                            // xcvr_native_s10_0:tx_clkout -> xcvr_st_converter_0:tx_clkout
	wire   [0:0] xcvr_native_s10_0_tx_clkout2_clk;                                                           // xcvr_native_s10_0:tx_clkout2 -> xcvr_test_system_0:xcvr_tx_rx_clkout2_converter_0_tx_clkout2_clk
	wire         xcvr_st_converter_0_tx_clkout_a_output_clk;                                                 // xcvr_st_converter_0:tx_clkout_a_output -> xcvr_native_s10_0:tx_coreclkin
	wire   [0:0] pll_locked_pll_locked_output_pll_locked;                                                    // pll_locked:pll_locked_output -> nativePHY_loopback_cont_0:pll_locked
	wire   [0:0] pll_locked_pll_locked_a_pll_locked;                                                         // pll_locked:pll_locked_a -> xcvr_reset_control_s10_0:pll_locked
	wire   [0:0] xcvr_reset_control_s10_0_rx_analogreset_rx_analogreset;                                     // xcvr_reset_control_s10_0:rx_analogreset -> xcvr_native_s10_0:rx_analogreset
	wire   [0:0] xcvr_native_s10_0_rx_analogreset_stat_rx_analogreset_stat;                                  // xcvr_native_s10_0:rx_analogreset_stat -> xcvr_reset_control_s10_0:rx_analogreset_stat
	wire   [0:0] xcvr_native_s10_0_rx_cal_busy_rx_cal_busy;                                                  // xcvr_native_s10_0:rx_cal_busy -> xcvr_reset_control_s10_0:rx_cal_busy
	wire         xcvr_st_converter_0_rx_clkout_a_export;                                                     // xcvr_st_converter_0:rx_clkout_a -> xcvr_test_system_0:xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_clk_export
	wire   [0:0] xcvr_reset_control_s10_0_rx_digitalreset_rx_digitalreset;                                   // xcvr_reset_control_s10_0:rx_digitalreset -> xcvr_native_s10_0:rx_digitalreset
	wire   [0:0] xcvr_native_s10_0_rx_digitalreset_stat_rx_digitalreset_stat;                                // xcvr_native_s10_0:rx_digitalreset_stat -> xcvr_reset_control_s10_0:rx_digitalreset_stat
	wire   [0:0] xcvr_native_s10_0_rx_is_lockedtodata_rx_is_lockedtodata;                                    // xcvr_native_s10_0:rx_is_lockedtodata -> xcvr_reset_control_s10_0:rx_is_lockedtodata
	wire   [0:0] xcvr_native_s10_0_rx_is_lockedtoref_rx_is_lockedtoref;                                      // xcvr_native_s10_0:rx_is_lockedtoref -> nativePHY_loopback_cont_0:rx_is_lockedtoref
	wire  [63:0] xcvr_native_s10_0_rx_parallel_data_rx_parallel_data;                                        // xcvr_native_s10_0:rx_parallel_data -> xcvr_st_converter_0:rx_parallel_data
	wire   [0:0] nativephy_loopback_cont_0_rx_seriallpbken_rx_seriallpbken;                                  // nativePHY_loopback_cont_0:rx_seriallpbken -> xcvr_native_s10_0:rx_seriallpbken
	wire   [0:0] xcvr_reset_control_s10_0_tx_analogreset_tx_analogreset;                                     // xcvr_reset_control_s10_0:tx_analogreset -> xcvr_native_s10_0:tx_analogreset
	wire   [0:0] xcvr_native_s10_0_tx_analogreset_stat_tx_analogreset_stat;                                  // xcvr_native_s10_0:tx_analogreset_stat -> xcvr_reset_control_s10_0:tx_analogreset_stat
	wire   [0:0] xcvr_native_s10_0_tx_cal_busy_tx_cal_busy;                                                  // xcvr_native_s10_0:tx_cal_busy -> xcvr_reset_control_s10_0:tx_cal_busy
	wire         xcvr_st_converter_0_tx_clkout_a_export;                                                     // xcvr_st_converter_0:tx_clkout_a -> xcvr_test_system_0:xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_clk_export
	wire   [0:0] xcvr_reset_control_s10_0_tx_digitalreset_tx_digitalreset;                                   // xcvr_reset_control_s10_0:tx_digitalreset -> xcvr_native_s10_0:tx_digitalreset
	wire   [0:0] xcvr_native_s10_0_tx_digitalreset_stat_tx_digitalreset_stat;                                // xcvr_native_s10_0:tx_digitalreset_stat -> xcvr_reset_control_s10_0:tx_digitalreset_stat
	wire  [63:0] xcvr_st_converter_0_tx_parallel_data_tx_parallel_data;                                      // xcvr_st_converter_0:tx_parallel_data -> xcvr_native_s10_0:tx_parallel_data
	wire  [63:0] xcvr_st_converter_0_rx_data_a_export;                                                       // xcvr_st_converter_0:rx_data_a -> xcvr_test_system_0:xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_export
	wire  [63:0] xcvr_test_system_0_xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_export; // xcvr_test_system_0:xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_export -> xcvr_st_converter_0:tx_data_a
	wire         clk_100_clk_reset_reset;                                                                    // clk_100:reset_n_out -> [rst_controller_001:reset_in0, xcvr_reset_control_s10_0:reset]
	wire         clk_50_clk_reset_reset;                                                                     // clk_50:reset_n_out -> [rst_controller:reset_in0, xcvr_test_system_0:reset_50_reset_n]
	wire  [31:0] default_pma_settings_conf_0_avalon_master_readdata;                                         // mm_interconnect_0:default_pma_settings_conf_0_avalon_master_readdata -> default_pma_settings_conf_0:master_rdata
	wire         default_pma_settings_conf_0_avalon_master_waitrequest;                                      // mm_interconnect_0:default_pma_settings_conf_0_avalon_master_waitrequest -> default_pma_settings_conf_0:waitrequest_in
	wire         default_pma_settings_conf_0_avalon_master_read;                                             // default_pma_settings_conf_0:master_oen -> mm_interconnect_0:default_pma_settings_conf_0_avalon_master_read
	wire   [3:0] default_pma_settings_conf_0_avalon_master_byteenable;                                       // default_pma_settings_conf_0:master_be -> mm_interconnect_0:default_pma_settings_conf_0_avalon_master_byteenable
	wire  [31:0] default_pma_settings_conf_0_avalon_master_address;                                          // default_pma_settings_conf_0:master_address -> mm_interconnect_0:default_pma_settings_conf_0_avalon_master_address
	wire         default_pma_settings_conf_0_avalon_master_readdatavalid;                                    // mm_interconnect_0:default_pma_settings_conf_0_avalon_master_readdatavalid -> default_pma_settings_conf_0:readdatavalid_in
	wire         default_pma_settings_conf_0_avalon_master_write;                                            // default_pma_settings_conf_0:master_wen -> mm_interconnect_0:default_pma_settings_conf_0_avalon_master_write
	wire  [31:0] default_pma_settings_conf_0_avalon_master_writedata;                                        // default_pma_settings_conf_0:master_wdata -> mm_interconnect_0:default_pma_settings_conf_0_avalon_master_writedata
	wire         mm_bridge_0_m0_waitrequest;                                                                 // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [31:0] mm_bridge_0_m0_readdata;                                                                    // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                                                 // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire  [14:0] mm_bridge_0_m0_address;                                                                     // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire         mm_bridge_0_m0_read;                                                                        // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire   [3:0] mm_bridge_0_m0_byteenable;                                                                  // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                                                               // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire  [31:0] mm_bridge_0_m0_writedata;                                                                   // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                                                       // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire   [0:0] mm_bridge_0_m0_burstcount;                                                                  // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire  [31:0] mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_readdata;                                 // xcvr_native_s10_0:reconfig_readdata -> mm_interconnect_0:xcvr_native_s10_0_reconfig_avmm_readdata
	wire         mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_waitrequest;                              // xcvr_native_s10_0:reconfig_waitrequest -> mm_interconnect_0:xcvr_native_s10_0_reconfig_avmm_waitrequest
	wire  [10:0] mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_address;                                  // mm_interconnect_0:xcvr_native_s10_0_reconfig_avmm_address -> xcvr_native_s10_0:reconfig_address
	wire         mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_read;                                     // mm_interconnect_0:xcvr_native_s10_0_reconfig_avmm_read -> xcvr_native_s10_0:reconfig_read
	wire         mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_write;                                    // mm_interconnect_0:xcvr_native_s10_0_reconfig_avmm_write -> xcvr_native_s10_0:reconfig_write
	wire  [31:0] mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_writedata;                                // mm_interconnect_0:xcvr_native_s10_0_reconfig_avmm_writedata -> xcvr_native_s10_0:reconfig_writedata
	wire  [31:0] mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_readdata;                        // default_pma_settings_conf_0:slave_readdata -> mm_interconnect_0:default_pma_settings_conf_0_avalon_slave_readdata
	wire   [3:0] mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_address;                         // mm_interconnect_0:default_pma_settings_conf_0_avalon_slave_address -> default_pma_settings_conf_0:slave_address
	wire         mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_read;                            // mm_interconnect_0:default_pma_settings_conf_0_avalon_slave_read -> default_pma_settings_conf_0:slave_read
	wire         mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_write;                           // mm_interconnect_0:default_pma_settings_conf_0_avalon_slave_write -> default_pma_settings_conf_0:slave_write
	wire  [31:0] mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_writedata;                       // mm_interconnect_0:default_pma_settings_conf_0_avalon_slave_writedata -> default_pma_settings_conf_0:slave_writedata
	wire  [31:0] mm_interconnect_0_nativephy_loopback_cont_0_csr_readdata;                                   // nativePHY_loopback_cont_0:csr_readdata -> mm_interconnect_0:nativePHY_loopback_cont_0_csr_readdata
	wire   [3:0] mm_interconnect_0_nativephy_loopback_cont_0_csr_address;                                    // mm_interconnect_0:nativePHY_loopback_cont_0_csr_address -> nativePHY_loopback_cont_0:csr_address
	wire         mm_interconnect_0_nativephy_loopback_cont_0_csr_read;                                       // mm_interconnect_0:nativePHY_loopback_cont_0_csr_read -> nativePHY_loopback_cont_0:csr_read
	wire         mm_interconnect_0_nativephy_loopback_cont_0_csr_write;                                      // mm_interconnect_0:nativePHY_loopback_cont_0_csr_write -> nativePHY_loopback_cont_0:csr_write
	wire  [31:0] mm_interconnect_0_nativephy_loopback_cont_0_csr_writedata;                                  // mm_interconnect_0:nativePHY_loopback_cont_0_csr_writedata -> nativePHY_loopback_cont_0:csr_writedata
	wire  [31:0] mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_readdata;                               // xcvr_test_system_0:mm_bridge_0_s0_readdata -> mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_waitrequest;                            // xcvr_test_system_0:mm_bridge_0_s0_waitrequest -> mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_waitrequest
	wire         mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_debugaccess;                            // mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_debugaccess -> xcvr_test_system_0:mm_bridge_0_s0_debugaccess
	wire  [12:0] mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_address;                                // mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_address -> xcvr_test_system_0:mm_bridge_0_s0_address
	wire         mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_read;                                   // mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_read -> xcvr_test_system_0:mm_bridge_0_s0_read
	wire   [3:0] mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_byteenable;                             // mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_byteenable -> xcvr_test_system_0:mm_bridge_0_s0_byteenable
	wire         mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_readdatavalid;                          // xcvr_test_system_0:mm_bridge_0_s0_readdatavalid -> mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_readdatavalid
	wire         mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_write;                                  // mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_write -> xcvr_test_system_0:mm_bridge_0_s0_write
	wire  [31:0] mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_writedata;                              // mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_writedata -> xcvr_test_system_0:mm_bridge_0_s0_writedata
	wire   [0:0] mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_burstcount;                             // mm_interconnect_0:xcvr_test_system_0_mm_bridge_0_s0_burstcount -> xcvr_test_system_0:mm_bridge_0_s0_burstcount
	wire         rst_controller_reset_out_reset;                                                             // rst_controller:reset_out -> [default_pma_settings_conf_0:reset_n, mm_bridge_0:reset, mm_interconnect_0:default_pma_settings_conf_0_reset_reset_bridge_in_reset_reset, nativePHY_loopback_cont_0:reset_n]
	wire         rst_controller_001_reset_out_reset;                                                         // rst_controller_001:reset_out -> [mm_interconnect_0:xcvr_native_s10_0_reconfig_reset_reset_bridge_in_reset_reset, xcvr_native_s10_0:reconfig_reset]

	qsfp_xcvr_test_clk_100 clk_100 (
		.in_clk      (clk_100_clk),             //   input,  width = 1,       clk_in.clk
		.reset_n     (reset_100_reset_n),       //   input,  width = 1, clk_in_reset.reset_n
		.clk_out     (clk_100_clk_clk),         //  output,  width = 1,          clk.clk
		.reset_n_out (clk_100_clk_reset_reset)  //  output,  width = 1,    clk_reset.reset_n
	);

	qsfp_xcvr_test_clk_50 clk_50 (
		.in_clk      (clk_50_clk),             //   input,  width = 1,       clk_in.clk
		.reset_n     (reset_50_reset_n),       //   input,  width = 1, clk_in_reset.reset_n
		.clk_out     (clk_50_clk_clk),         //  output,  width = 1,          clk.clk
		.reset_n_out (clk_50_clk_reset_reset)  //  output,  width = 1,    clk_reset.reset_n
	);

	qsfp_xcvr_test_default_pma_settings_conf_0 default_pma_settings_conf_0 (
		.clock            (clk_50_clk_clk),                                                       //   input,   width = 1,         clock.clk
		.reset_n          (~rst_controller_reset_out_reset),                                      //   input,   width = 1,         reset.reset_n
		.master_wen       (default_pma_settings_conf_0_avalon_master_write),                      //  output,   width = 1, avalon_master.write_n
		.master_oen       (default_pma_settings_conf_0_avalon_master_read),                       //  output,   width = 1,              .read_n
		.master_be        (default_pma_settings_conf_0_avalon_master_byteenable),                 //  output,   width = 4,              .byteenable
		.master_address   (default_pma_settings_conf_0_avalon_master_address),                    //  output,  width = 32,              .address
		.master_wdata     (default_pma_settings_conf_0_avalon_master_writedata),                  //  output,  width = 32,              .writedata
		.master_rdata     (default_pma_settings_conf_0_avalon_master_readdata),                   //   input,  width = 32,              .readdata
		.readdatavalid_in (default_pma_settings_conf_0_avalon_master_readdatavalid),              //   input,   width = 1,              .readdatavalid
		.waitrequest_in   (default_pma_settings_conf_0_avalon_master_waitrequest),                //   input,   width = 1,              .waitrequest
		.slave_read       (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_read),      //   input,   width = 1,  avalon_slave.read
		.slave_write      (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_write),     //   input,   width = 1,              .write
		.slave_readdata   (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_readdata),  //  output,  width = 32,              .readdata
		.slave_writedata  (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_writedata), //   input,  width = 32,              .writedata
		.slave_address    (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_address)    //   input,   width = 4,              .address
	);

	qsfp_xcvr_test_mm_bridge_0 mm_bridge_0 (
		.clk              (clk_50_clk_clk),                 //   input,   width = 1,   clk.clk
		.reset            (rst_controller_reset_out_reset), //   input,   width = 1, reset.reset
		.s0_waitrequest   (mm_bridge_0_s0_waitrequest),     //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (mm_bridge_0_s0_readdata),        //  output,  width = 32,      .readdata
		.s0_readdatavalid (mm_bridge_0_s0_readdatavalid),   //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (mm_bridge_0_s0_burstcount),      //   input,   width = 1,      .burstcount
		.s0_writedata     (mm_bridge_0_s0_writedata),       //   input,  width = 32,      .writedata
		.s0_address       (mm_bridge_0_s0_address),         //   input,  width = 15,      .address
		.s0_write         (mm_bridge_0_s0_write),           //   input,   width = 1,      .write
		.s0_read          (mm_bridge_0_s0_read),            //   input,   width = 1,      .read
		.s0_byteenable    (mm_bridge_0_s0_byteenable),      //   input,   width = 4,      .byteenable
		.s0_debugaccess   (mm_bridge_0_s0_debugaccess),     //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),        //   input,  width = 32,      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),      //  output,   width = 1,      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),       //  output,  width = 32,      .writedata
		.m0_address       (mm_bridge_0_m0_address),         //  output,  width = 15,      .address
		.m0_write         (mm_bridge_0_m0_write),           //  output,   width = 1,      .write
		.m0_read          (mm_bridge_0_m0_read),            //  output,   width = 1,      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),      //  output,   width = 4,      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess)      //  output,   width = 1,      .debugaccess
	);

	qsfp_xcvr_test_nativePHY_loopback_cont_0 nativephy_loopback_cont_0 (
		.reset_n             (~rst_controller_reset_out_reset),                           //   input,   width = 1,               reset.reset_n
		.clk                 (clk_50_clk_clk),                                            //   input,   width = 1,               clock.clk
		.csr_address         (mm_interconnect_0_nativephy_loopback_cont_0_csr_address),   //   input,   width = 4,                 csr.address
		.csr_read            (mm_interconnect_0_nativephy_loopback_cont_0_csr_read),      //   input,   width = 1,                    .read
		.csr_write           (mm_interconnect_0_nativephy_loopback_cont_0_csr_write),     //   input,   width = 1,                    .write
		.csr_readdata        (mm_interconnect_0_nativephy_loopback_cont_0_csr_readdata),  //  output,  width = 32,                    .readdata
		.csr_writedata       (mm_interconnect_0_nativephy_loopback_cont_0_csr_writedata), //   input,  width = 32,                    .writedata
		.pll_locked          (pll_locked_pll_locked_output_pll_locked),                   //   input,   width = 1,          pll_locked.pll_locked
		.rx_is_lockedtoref   (xcvr_native_s10_0_rx_is_lockedtoref_rx_is_lockedtoref),     //   input,   width = 1,   rx_is_lockedtoref.rx_is_lockedtoref
		.rx_seriallpbken     (nativephy_loopback_cont_0_rx_seriallpbken_rx_seriallpbken), //  output,   width = 1,     rx_seriallpbken.rx_seriallpbken
		.rx_seriallpbken_mon ()                                                           //  output,   width = 1, rx_seriallpbken_mon.export
	);

	qsfp_xcvr_test_pll_status_interconnect_0 pll_locked (
		.pll_locked        (pll_locked_pll_locked_pll_locked),        //   input,  width = 1,        pll_locked.pll_locked
		.pll_powerdown     (),                                        //  output,  width = 1,     pll_powerdown.pll_powerdown
		.mcgb_rst          (),                                        //  output,  width = 1,          mcgb_rst.mcgb_rst
		.pll_locked_output (pll_locked_pll_locked_output_pll_locked), //  output,  width = 1, pll_locked_output.pll_locked
		.pll_locked_a      (pll_locked_pll_locked_a_pll_locked),      //  output,  width = 1,      pll_locked_a.pll_locked
		.pll_powerdown_a   ()                                         //   input,  width = 1,   pll_powerdown_a.pll_powerdown
	);

	qsfp_xcvr_test_xcvr_native_s10_htile_1 xcvr_native_s10_0 (
		.tx_analogreset          (xcvr_reset_control_s10_0_tx_analogreset_tx_analogreset),        //   input,   width = 1,          tx_analogreset.tx_analogreset
		.rx_analogreset          (xcvr_reset_control_s10_0_rx_analogreset_rx_analogreset),        //   input,   width = 1,          rx_analogreset.rx_analogreset
		.tx_digitalreset         (xcvr_reset_control_s10_0_tx_digitalreset_tx_digitalreset),      //   input,   width = 1,         tx_digitalreset.tx_digitalreset
		.rx_digitalreset         (xcvr_reset_control_s10_0_rx_digitalreset_rx_digitalreset),      //   input,   width = 1,         rx_digitalreset.rx_digitalreset
		.tx_analogreset_stat     (xcvr_native_s10_0_tx_analogreset_stat_tx_analogreset_stat),     //  output,   width = 1,     tx_analogreset_stat.tx_analogreset_stat
		.rx_analogreset_stat     (xcvr_native_s10_0_rx_analogreset_stat_rx_analogreset_stat),     //  output,   width = 1,     rx_analogreset_stat.rx_analogreset_stat
		.tx_digitalreset_stat    (xcvr_native_s10_0_tx_digitalreset_stat_tx_digitalreset_stat),   //  output,   width = 1,    tx_digitalreset_stat.tx_digitalreset_stat
		.rx_digitalreset_stat    (xcvr_native_s10_0_rx_digitalreset_stat_rx_digitalreset_stat),   //  output,   width = 1,    rx_digitalreset_stat.rx_digitalreset_stat
		.tx_cal_busy             (xcvr_native_s10_0_tx_cal_busy_tx_cal_busy),                     //  output,   width = 1,             tx_cal_busy.tx_cal_busy
		.rx_cal_busy             (xcvr_native_s10_0_rx_cal_busy_rx_cal_busy),                     //  output,   width = 1,             rx_cal_busy.rx_cal_busy
		.tx_serial_clk0          (xcvr_native_s10_0_tx_serial_clk0_clk),                          //   input,   width = 1,          tx_serial_clk0.clk
		.rx_cdr_refclk0          (xcvr_native_s10_0_rx_cdr_refclk0_clk),                          //   input,   width = 1,          rx_cdr_refclk0.clk
		.tx_serial_data          (xcvr_native_s10_0_tx_serial_data_tx_serial_data),               //  output,   width = 1,          tx_serial_data.tx_serial_data
		.rx_serial_data          (xcvr_native_s10_0_rx_serial_data_rx_serial_data),               //   input,   width = 1,          rx_serial_data.rx_serial_data
		.rx_seriallpbken         (nativephy_loopback_cont_0_rx_seriallpbken_rx_seriallpbken),     //   input,   width = 1,         rx_seriallpbken.rx_seriallpbken
		.rx_is_lockedtoref       (xcvr_native_s10_0_rx_is_lockedtoref_rx_is_lockedtoref),         //  output,   width = 1,       rx_is_lockedtoref.rx_is_lockedtoref
		.rx_is_lockedtodata      (xcvr_native_s10_0_rx_is_lockedtodata_rx_is_lockedtodata),       //  output,   width = 1,      rx_is_lockedtodata.rx_is_lockedtodata
		.tx_coreclkin            (xcvr_st_converter_0_tx_clkout_a_output_clk),                    //   input,   width = 1,            tx_coreclkin.clk
		.rx_coreclkin            (xcvr_st_converter_0_rx_clkout_a_output_clk),                    //   input,   width = 1,            rx_coreclkin.clk
		.tx_clkout               (xcvr_native_s10_0_tx_clkout_clk),                               //  output,   width = 1,               tx_clkout.clk
		.tx_clkout2              (xcvr_native_s10_0_tx_clkout2_clk),                              //  output,   width = 1,              tx_clkout2.clk
		.rx_clkout               (xcvr_native_s10_0_rx_clkout_clk),                               //  output,   width = 1,               rx_clkout.clk
		.rx_clkout2              (xcvr_native_s10_0_rx_clkout2_clk),                              //  output,   width = 1,              rx_clkout2.clk
		.rx_pma_iqtxrx_clkout    (),                                                              //  output,   width = 1,    rx_pma_iqtxrx_clkout.clk
		.tx_parallel_data        (xcvr_st_converter_0_tx_parallel_data_tx_parallel_data),         //   input,  width = 64,        tx_parallel_data.tx_parallel_data
		.unused_tx_parallel_data (),                                                              //   input,  width = 16, unused_tx_parallel_data.unused_tx_parallel_data
		.rx_parallel_data        (xcvr_native_s10_0_rx_parallel_data_rx_parallel_data),           //  output,  width = 64,        rx_parallel_data.rx_parallel_data
		.unused_rx_parallel_data (),                                                              //  output,  width = 16, unused_rx_parallel_data.unused_rx_parallel_data
		.reconfig_clk            (clk_100_clk_clk),                                               //   input,   width = 1,            reconfig_clk.clk
		.reconfig_reset          (rst_controller_001_reset_out_reset),                            //   input,   width = 1,          reconfig_reset.reset
		.reconfig_write          (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_write),       //   input,   width = 1,           reconfig_avmm.write
		.reconfig_read           (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_read),        //   input,   width = 1,                        .read
		.reconfig_address        (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_address),     //   input,  width = 11,                        .address
		.reconfig_writedata      (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_writedata),   //   input,  width = 32,                        .writedata
		.reconfig_readdata       (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_readdata),    //  output,  width = 32,                        .readdata
		.reconfig_waitrequest    (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_waitrequest)  //  output,   width = 1,                        .waitrequest
	);

	qsfp_xcvr_test_xcvr_reset_control_s10_0 xcvr_reset_control_s10_0 (
		.clock                (clk_100_clk_clk),                                             //   input,  width = 1,                clock.clk
		.reset                (~clk_100_clk_reset_reset),                                    //   input,  width = 1,                reset.reset
		.tx_analogreset       (xcvr_reset_control_s10_0_tx_analogreset_tx_analogreset),      //  output,  width = 1,       tx_analogreset.tx_analogreset
		.tx_digitalreset      (xcvr_reset_control_s10_0_tx_digitalreset_tx_digitalreset),    //  output,  width = 1,      tx_digitalreset.tx_digitalreset
		.tx_ready             (),                                                            //  output,  width = 1,             tx_ready.tx_ready
		.pll_locked           (pll_locked_pll_locked_a_pll_locked),                          //   input,  width = 1,           pll_locked.pll_locked
		.pll_select           (),                                                            //   input,  width = 1,           pll_select.pll_select
		.tx_cal_busy          (xcvr_native_s10_0_tx_cal_busy_tx_cal_busy),                   //   input,  width = 1,          tx_cal_busy.tx_cal_busy
		.tx_analogreset_stat  (xcvr_native_s10_0_tx_analogreset_stat_tx_analogreset_stat),   //   input,  width = 1,  tx_analogreset_stat.tx_analogreset_stat
		.tx_digitalreset_stat (xcvr_native_s10_0_tx_digitalreset_stat_tx_digitalreset_stat), //   input,  width = 1, tx_digitalreset_stat.tx_digitalreset_stat
		.rx_analogreset       (xcvr_reset_control_s10_0_rx_analogreset_rx_analogreset),      //  output,  width = 1,       rx_analogreset.rx_analogreset
		.rx_digitalreset      (xcvr_reset_control_s10_0_rx_digitalreset_rx_digitalreset),    //  output,  width = 1,      rx_digitalreset.rx_digitalreset
		.rx_ready             (),                                                            //  output,  width = 1,             rx_ready.rx_ready
		.rx_is_lockedtodata   (xcvr_native_s10_0_rx_is_lockedtodata_rx_is_lockedtodata),     //   input,  width = 1,   rx_is_lockedtodata.rx_is_lockedtodata
		.rx_cal_busy          (xcvr_native_s10_0_rx_cal_busy_rx_cal_busy),                   //   input,  width = 1,          rx_cal_busy.rx_cal_busy
		.rx_analogreset_stat  (xcvr_native_s10_0_rx_analogreset_stat_rx_analogreset_stat),   //   input,  width = 1,  rx_analogreset_stat.rx_analogreset_stat
		.rx_digitalreset_stat (xcvr_native_s10_0_rx_digitalreset_stat_rx_digitalreset_stat)  //   input,  width = 1, rx_digitalreset_stat.rx_digitalreset_stat
	);

	qsfp_xcvr_test_xcvr_st_converter_0 xcvr_st_converter_0 (
		.tx_parallel_data   (xcvr_st_converter_0_tx_parallel_data_tx_parallel_data),                                      //  output,  width = 64,   tx_parallel_data.tx_parallel_data
		.tx_clkout          (xcvr_native_s10_0_tx_clkout_clk),                                                            //   input,   width = 1,          tx_clkout.clk
		.rx_parallel_data   (xcvr_native_s10_0_rx_parallel_data_rx_parallel_data),                                        //   input,  width = 64,   rx_parallel_data.rx_parallel_data
		.rx_clkout          (xcvr_native_s10_0_rx_clkout_clk),                                                            //   input,   width = 1,          rx_clkout.clk
		.rx_is_lockedtodata (),                                                                                           //   input,   width = 1, rx_is_lockedtodata.rx_is_lockedtodata
		.tx_data_a          (xcvr_test_system_0_xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_export), //   input,  width = 64,          tx_data_a.export
		.tx_clkout_a        (xcvr_st_converter_0_tx_clkout_a_export),                                                     //  output,   width = 1,        tx_clkout_a.export
		.rx_data_a          (xcvr_st_converter_0_rx_data_a_export),                                                       //  output,  width = 64,          rx_data_a.export
		.rx_clkout_a        (xcvr_st_converter_0_rx_clkout_a_export),                                                     //  output,   width = 1,        rx_clkout_a.export
		.test_reset_n_a     (),                                                                                           //  output,   width = 1,     test_reset_n_a.reset_n
		.tx_clkout_a_output (xcvr_st_converter_0_tx_clkout_a_output_clk),                                                 //  output,   width = 1, tx_clkout_a_output.clk
		.rx_clkout_a_output (xcvr_st_converter_0_rx_clkout_a_output_clk)                                                  //  output,   width = 1, rx_clkout_a_output.clk
	);

	xcvr_test_system xcvr_test_system_0 (
		.clk_50_clk                                                                  (clk_50_clk_clk),                                                                             //   input,   width = 1,                                                               clk_50.clk
		.reset_50_reset_n                                                            (clk_50_clk_reset_reset),                                                                     //   input,   width = 1,                                                             reset_50.reset_n
		.mm_bridge_0_s0_waitrequest                                                  (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_waitrequest),                            //  output,   width = 1,                                                       mm_bridge_0_s0.waitrequest
		.mm_bridge_0_s0_readdata                                                     (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_readdata),                               //  output,  width = 32,                                                                     .readdata
		.mm_bridge_0_s0_readdatavalid                                                (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_readdatavalid),                          //  output,   width = 1,                                                                     .readdatavalid
		.mm_bridge_0_s0_burstcount                                                   (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_burstcount),                             //   input,   width = 1,                                                                     .burstcount
		.mm_bridge_0_s0_writedata                                                    (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_writedata),                              //   input,  width = 32,                                                                     .writedata
		.mm_bridge_0_s0_address                                                      (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_address),                                //   input,  width = 13,                                                                     .address
		.mm_bridge_0_s0_write                                                        (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_write),                                  //   input,   width = 1,                                                                     .write
		.mm_bridge_0_s0_read                                                         (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_read),                                   //   input,   width = 1,                                                                     .read
		.mm_bridge_0_s0_byteenable                                                   (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_byteenable),                             //   input,   width = 4,                                                                     .byteenable
		.mm_bridge_0_s0_debugaccess                                                  (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_debugaccess),                            //   input,   width = 1,                                                                     .debugaccess
		.xcvr_tx_rx_clkout2_converter_0_rx_clkout2_clk                               (xcvr_native_s10_0_rx_clkout2_clk),                                                           //   input,   width = 1,                            xcvr_tx_rx_clkout2_converter_0_rx_clkout2.clk
		.xcvr_tx_rx_clkout2_converter_0_tx_clkout2_clk                               (xcvr_native_s10_0_tx_clkout2_clk),                                                           //   input,   width = 1,                            xcvr_tx_rx_clkout2_converter_0_tx_clkout2.clk
		.xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_export        (xcvr_st_converter_0_rx_data_a_export),                                                       //   input,  width = 64,        xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in.export
		.xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_clk_export    (xcvr_st_converter_0_rx_clkout_a_export),                                                     //   input,   width = 1,    xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_clk.export
		.xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_export     (xcvr_test_system_0_xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_export), //  output,  width = 64,     xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out.export
		.xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_clk_export (xcvr_st_converter_0_tx_clkout_a_export)                                                      //   input,   width = 1, xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_clk.export
	);

	qsfp_xcvr_test_altera_mm_interconnect_1920_4ix6v3i mm_interconnect_0 (
		.default_pma_settings_conf_0_avalon_master_address             (default_pma_settings_conf_0_avalon_master_address),                    //   input,  width = 32,               default_pma_settings_conf_0_avalon_master.address
		.default_pma_settings_conf_0_avalon_master_waitrequest         (default_pma_settings_conf_0_avalon_master_waitrequest),                //  output,   width = 1,                                                        .waitrequest
		.default_pma_settings_conf_0_avalon_master_byteenable          (default_pma_settings_conf_0_avalon_master_byteenable),                 //   input,   width = 4,                                                        .byteenable
		.default_pma_settings_conf_0_avalon_master_read                (~default_pma_settings_conf_0_avalon_master_read),                      //   input,   width = 1,                                                        .read
		.default_pma_settings_conf_0_avalon_master_readdata            (default_pma_settings_conf_0_avalon_master_readdata),                   //  output,  width = 32,                                                        .readdata
		.default_pma_settings_conf_0_avalon_master_readdatavalid       (default_pma_settings_conf_0_avalon_master_readdatavalid),              //  output,   width = 1,                                                        .readdatavalid
		.default_pma_settings_conf_0_avalon_master_write               (~default_pma_settings_conf_0_avalon_master_write),                     //   input,   width = 1,                                                        .write
		.default_pma_settings_conf_0_avalon_master_writedata           (default_pma_settings_conf_0_avalon_master_writedata),                  //   input,  width = 32,                                                        .writedata
		.mm_bridge_0_m0_address                                        (mm_bridge_0_m0_address),                                               //   input,  width = 15,                                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                                    (mm_bridge_0_m0_waitrequest),                                           //  output,   width = 1,                                                        .waitrequest
		.mm_bridge_0_m0_burstcount                                     (mm_bridge_0_m0_burstcount),                                            //   input,   width = 1,                                                        .burstcount
		.mm_bridge_0_m0_byteenable                                     (mm_bridge_0_m0_byteenable),                                            //   input,   width = 4,                                                        .byteenable
		.mm_bridge_0_m0_read                                           (mm_bridge_0_m0_read),                                                  //   input,   width = 1,                                                        .read
		.mm_bridge_0_m0_readdata                                       (mm_bridge_0_m0_readdata),                                              //  output,  width = 32,                                                        .readdata
		.mm_bridge_0_m0_readdatavalid                                  (mm_bridge_0_m0_readdatavalid),                                         //  output,   width = 1,                                                        .readdatavalid
		.mm_bridge_0_m0_write                                          (mm_bridge_0_m0_write),                                                 //   input,   width = 1,                                                        .write
		.mm_bridge_0_m0_writedata                                      (mm_bridge_0_m0_writedata),                                             //   input,  width = 32,                                                        .writedata
		.mm_bridge_0_m0_debugaccess                                    (mm_bridge_0_m0_debugaccess),                                           //   input,   width = 1,                                                        .debugaccess
		.xcvr_native_s10_0_reconfig_avmm_address                       (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_address),            //  output,  width = 11,                         xcvr_native_s10_0_reconfig_avmm.address
		.xcvr_native_s10_0_reconfig_avmm_write                         (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_write),              //  output,   width = 1,                                                        .write
		.xcvr_native_s10_0_reconfig_avmm_read                          (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_read),               //  output,   width = 1,                                                        .read
		.xcvr_native_s10_0_reconfig_avmm_readdata                      (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_readdata),           //   input,  width = 32,                                                        .readdata
		.xcvr_native_s10_0_reconfig_avmm_writedata                     (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_writedata),          //  output,  width = 32,                                                        .writedata
		.xcvr_native_s10_0_reconfig_avmm_waitrequest                   (mm_interconnect_0_xcvr_native_s10_0_reconfig_avmm_waitrequest),        //   input,   width = 1,                                                        .waitrequest
		.default_pma_settings_conf_0_avalon_slave_address              (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_address),   //  output,   width = 4,                default_pma_settings_conf_0_avalon_slave.address
		.default_pma_settings_conf_0_avalon_slave_write                (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_write),     //  output,   width = 1,                                                        .write
		.default_pma_settings_conf_0_avalon_slave_read                 (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_read),      //  output,   width = 1,                                                        .read
		.default_pma_settings_conf_0_avalon_slave_readdata             (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_readdata),  //   input,  width = 32,                                                        .readdata
		.default_pma_settings_conf_0_avalon_slave_writedata            (mm_interconnect_0_default_pma_settings_conf_0_avalon_slave_writedata), //  output,  width = 32,                                                        .writedata
		.nativePHY_loopback_cont_0_csr_address                         (mm_interconnect_0_nativephy_loopback_cont_0_csr_address),              //  output,   width = 4,                           nativePHY_loopback_cont_0_csr.address
		.nativePHY_loopback_cont_0_csr_write                           (mm_interconnect_0_nativephy_loopback_cont_0_csr_write),                //  output,   width = 1,                                                        .write
		.nativePHY_loopback_cont_0_csr_read                            (mm_interconnect_0_nativephy_loopback_cont_0_csr_read),                 //  output,   width = 1,                                                        .read
		.nativePHY_loopback_cont_0_csr_readdata                        (mm_interconnect_0_nativephy_loopback_cont_0_csr_readdata),             //   input,  width = 32,                                                        .readdata
		.nativePHY_loopback_cont_0_csr_writedata                       (mm_interconnect_0_nativephy_loopback_cont_0_csr_writedata),            //  output,  width = 32,                                                        .writedata
		.xcvr_test_system_0_mm_bridge_0_s0_address                     (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_address),          //  output,  width = 13,                       xcvr_test_system_0_mm_bridge_0_s0.address
		.xcvr_test_system_0_mm_bridge_0_s0_write                       (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_write),            //  output,   width = 1,                                                        .write
		.xcvr_test_system_0_mm_bridge_0_s0_read                        (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_read),             //  output,   width = 1,                                                        .read
		.xcvr_test_system_0_mm_bridge_0_s0_readdata                    (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_readdata),         //   input,  width = 32,                                                        .readdata
		.xcvr_test_system_0_mm_bridge_0_s0_writedata                   (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_writedata),        //  output,  width = 32,                                                        .writedata
		.xcvr_test_system_0_mm_bridge_0_s0_burstcount                  (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_burstcount),       //  output,   width = 1,                                                        .burstcount
		.xcvr_test_system_0_mm_bridge_0_s0_byteenable                  (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_byteenable),       //  output,   width = 4,                                                        .byteenable
		.xcvr_test_system_0_mm_bridge_0_s0_readdatavalid               (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_readdatavalid),    //   input,   width = 1,                                                        .readdatavalid
		.xcvr_test_system_0_mm_bridge_0_s0_waitrequest                 (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_waitrequest),      //   input,   width = 1,                                                        .waitrequest
		.xcvr_test_system_0_mm_bridge_0_s0_debugaccess                 (mm_interconnect_0_xcvr_test_system_0_mm_bridge_0_s0_debugaccess),      //  output,   width = 1,                                                        .debugaccess
		.default_pma_settings_conf_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                       //   input,   width = 1, default_pma_settings_conf_0_reset_reset_bridge_in_reset.reset
		.xcvr_native_s10_0_reconfig_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                                   //   input,   width = 1,  xcvr_native_s10_0_reconfig_reset_reset_bridge_in_reset.reset
		.clk_50_clk_clk                                                (clk_50_clk_clk),                                                       //   input,   width = 1,                                              clk_50_clk.clk
		.clk_100_clk_clk                                               (clk_100_clk_clk)                                                       //   input,   width = 1,                                             clk_100_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clk_50_clk_reset_reset),        //   input,  width = 1, reset_in0.reset
		.clk            (clk_50_clk_clk),                 //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~clk_100_clk_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (clk_100_clk_clk),                    //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
