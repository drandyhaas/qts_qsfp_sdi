// xcvr_test_system.v

// Generated using ACDS version 23.3 104

`timescale 1 ps / 1 ps
module xcvr_test_system (
		input  wire        clk_50_clk,                                                                  //                                                               clk_50.clk
		input  wire        reset_50_reset_n,                                                            //                                                             reset_50.reset_n
		output wire        mm_bridge_0_s0_waitrequest,                                                  //                                                       mm_bridge_0_s0.waitrequest
		output wire [31:0] mm_bridge_0_s0_readdata,                                                     //                                                                     .readdata
		output wire        mm_bridge_0_s0_readdatavalid,                                                //                                                                     .readdatavalid
		input  wire [0:0]  mm_bridge_0_s0_burstcount,                                                   //                                                                     .burstcount
		input  wire [31:0] mm_bridge_0_s0_writedata,                                                    //                                                                     .writedata
		input  wire [12:0] mm_bridge_0_s0_address,                                                      //                                                                     .address
		input  wire        mm_bridge_0_s0_write,                                                        //                                                                     .write
		input  wire        mm_bridge_0_s0_read,                                                         //                                                                     .read
		input  wire [3:0]  mm_bridge_0_s0_byteenable,                                                   //                                                                     .byteenable
		input  wire        mm_bridge_0_s0_debugaccess,                                                  //                                                                     .debugaccess
		input  wire        xcvr_tx_rx_clkout2_converter_0_rx_clkout2_clk,                               //                            xcvr_tx_rx_clkout2_converter_0_rx_clkout2.clk
		input  wire        xcvr_tx_rx_clkout2_converter_0_tx_clkout2_clk,                               //                            xcvr_tx_rx_clkout2_converter_0_tx_clkout2.clk
		input  wire [63:0] xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_export,        //        xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in.export
		input  wire        xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_clk_export,    //    xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_clk.export
		output wire [63:0] xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_export,     //     xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out.export
		input  wire        xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_clk_export  // xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_clk.export
	);

	wire          clk_50_clk_clk;                                                                 // clk_50:clk_out -> [data_pattern_checker_0:csr_clk_clk, data_pattern_generator_0:csr_clk_clk, freq_counter_0:clk, mm_bridge_0:clk, mm_interconnect_0:clk_50_clk_clk, rst_controller:clk]
	wire          xcvr_tx_rx_clkout2_converter_0_tx_clkout2_sample_clk;                           // xcvr_tx_rx_clkout2_converter_0:tx_clkout2_sample -> freq_counter_0:sample_clk
	wire  [127:0] xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_fifo_read_export; // xcvr_user_rx_fifo_converter_0:data_pattern_checker_pattern_in_fifo_read -> data_pattern_checker_0:asi_data
	wire          xcvr_tx_rx_clkout2_converter_0_rx_clkout2_a_export;                             // xcvr_tx_rx_clkout2_converter_0:rx_clkout2_a -> data_pattern_checker_0:conduit_pattern_in_clk_export
	wire  [127:0] data_pattern_generator_0_conduit_pattern_out_export;                            // data_pattern_generator_0:aso_data -> xcvr_user_tx_fifo_converter_0:data_pattern_generator_pattern_out_fifo_write
	wire          xcvr_tx_rx_clkout2_converter_0_tx_clkout2_a_export;                             // xcvr_tx_rx_clkout2_converter_0:tx_clkout2_a -> data_pattern_generator_0:conduit_pattern_out_clk_export
	wire          xcvr_user_tx_fifo_converter_0_fifo_input_wrreq;                                 // xcvr_user_tx_fifo_converter_0:wrreq -> tx_fifo:wrreq
	wire          xcvr_user_tx_fifo_converter_0_fifo_input_wrclk;                                 // xcvr_user_tx_fifo_converter_0:wrclk -> tx_fifo:wrclk
	wire          xcvr_user_tx_fifo_converter_0_fifo_input_rdclk;                                 // xcvr_user_tx_fifo_converter_0:rdclk -> tx_fifo:rdclk
	wire          xcvr_user_tx_fifo_converter_0_fifo_input_rdreq;                                 // xcvr_user_tx_fifo_converter_0:rdreq -> tx_fifo:rdreq
	wire  [127:0] xcvr_user_tx_fifo_converter_0_fifo_input_datain;                                // xcvr_user_tx_fifo_converter_0:data -> tx_fifo:data
	wire          xcvr_user_rx_fifo_converter_0_fifo_input_wrreq;                                 // xcvr_user_rx_fifo_converter_0:wrreq -> rx_fifo:wrreq
	wire          xcvr_user_rx_fifo_converter_0_fifo_input_wrclk;                                 // xcvr_user_rx_fifo_converter_0:wrclk -> rx_fifo:wrclk
	wire          xcvr_user_rx_fifo_converter_0_fifo_input_rdclk;                                 // xcvr_user_rx_fifo_converter_0:rdclk -> rx_fifo:rdclk
	wire          xcvr_user_rx_fifo_converter_0_fifo_input_rdreq;                                 // xcvr_user_rx_fifo_converter_0:rdreq -> rx_fifo:rdreq
	wire   [63:0] xcvr_user_rx_fifo_converter_0_fifo_input_datain;                                // xcvr_user_rx_fifo_converter_0:data -> rx_fifo:data
	wire   [63:0] tx_fifo_fifo_output_dataout;                                                    // tx_fifo:q -> xcvr_user_tx_fifo_converter_0:q
	wire          tx_fifo_fifo_output_rdempty;                                                    // tx_fifo:rdempty -> xcvr_user_tx_fifo_converter_0:rdempty
	wire          tx_fifo_fifo_output_wrfull;                                                     // tx_fifo:wrfull -> xcvr_user_tx_fifo_converter_0:wrfull
	wire  [127:0] rx_fifo_fifo_output_dataout;                                                    // rx_fifo:q -> xcvr_user_rx_fifo_converter_0:q
	wire          rx_fifo_fifo_output_rdempty;                                                    // rx_fifo:rdempty -> xcvr_user_rx_fifo_converter_0:rdempty
	wire          rx_fifo_fifo_output_wrfull;                                                     // rx_fifo:wrfull -> xcvr_user_rx_fifo_converter_0:wrfull
	wire          xcvr_tx_rx_clkout2_converter_0_rx_clkout2_b_export;                             // xcvr_tx_rx_clkout2_converter_0:rx_clkout2_b -> xcvr_user_rx_fifo_converter_0:data_pattern_checker_pattern_in_fifo_read_clk
	wire          xcvr_tx_rx_clkout2_converter_0_tx_clkout2_b_export;                             // xcvr_tx_rx_clkout2_converter_0:tx_clkout2_b -> xcvr_user_tx_fifo_converter_0:data_pattern_generator_pattern_out_fifo_write_clk
	wire          mm_bridge_0_m0_waitrequest;                                                     // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire   [31:0] mm_bridge_0_m0_readdata;                                                        // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire          mm_bridge_0_m0_debugaccess;                                                     // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire   [12:0] mm_bridge_0_m0_address;                                                         // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire          mm_bridge_0_m0_read;                                                            // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire    [3:0] mm_bridge_0_m0_byteenable;                                                      // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire          mm_bridge_0_m0_readdatavalid;                                                   // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire   [31:0] mm_bridge_0_m0_writedata;                                                       // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire          mm_bridge_0_m0_write;                                                           // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire    [0:0] mm_bridge_0_m0_burstcount;                                                      // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire   [31:0] mm_interconnect_0_freq_counter_0_csr_readdata;                                  // freq_counter_0:csr_readdata -> mm_interconnect_0:freq_counter_0_csr_readdata
	wire    [3:0] mm_interconnect_0_freq_counter_0_csr_address;                                   // mm_interconnect_0:freq_counter_0_csr_address -> freq_counter_0:csr_address
	wire          mm_interconnect_0_freq_counter_0_csr_read;                                      // mm_interconnect_0:freq_counter_0_csr_read -> freq_counter_0:csr_read
	wire   [31:0] mm_interconnect_0_data_pattern_generator_0_csr_slave_readdata;                  // data_pattern_generator_0:csr_slave_readdata -> mm_interconnect_0:data_pattern_generator_0_csr_slave_readdata
	wire    [2:0] mm_interconnect_0_data_pattern_generator_0_csr_slave_address;                   // mm_interconnect_0:data_pattern_generator_0_csr_slave_address -> data_pattern_generator_0:csr_slave_address
	wire          mm_interconnect_0_data_pattern_generator_0_csr_slave_read;                      // mm_interconnect_0:data_pattern_generator_0_csr_slave_read -> data_pattern_generator_0:csr_slave_read
	wire    [3:0] mm_interconnect_0_data_pattern_generator_0_csr_slave_byteenable;                // mm_interconnect_0:data_pattern_generator_0_csr_slave_byteenable -> data_pattern_generator_0:csr_slave_byteenable
	wire          mm_interconnect_0_data_pattern_generator_0_csr_slave_write;                     // mm_interconnect_0:data_pattern_generator_0_csr_slave_write -> data_pattern_generator_0:csr_slave_write
	wire   [31:0] mm_interconnect_0_data_pattern_generator_0_csr_slave_writedata;                 // mm_interconnect_0:data_pattern_generator_0_csr_slave_writedata -> data_pattern_generator_0:csr_slave_writedata
	wire   [31:0] mm_interconnect_0_data_pattern_checker_0_csr_slave_readdata;                    // data_pattern_checker_0:csr_slave_readdata -> mm_interconnect_0:data_pattern_checker_0_csr_slave_readdata
	wire    [2:0] mm_interconnect_0_data_pattern_checker_0_csr_slave_address;                     // mm_interconnect_0:data_pattern_checker_0_csr_slave_address -> data_pattern_checker_0:csr_slave_address
	wire          mm_interconnect_0_data_pattern_checker_0_csr_slave_read;                        // mm_interconnect_0:data_pattern_checker_0_csr_slave_read -> data_pattern_checker_0:csr_slave_read
	wire    [3:0] mm_interconnect_0_data_pattern_checker_0_csr_slave_byteenable;                  // mm_interconnect_0:data_pattern_checker_0_csr_slave_byteenable -> data_pattern_checker_0:csr_slave_byteenable
	wire          mm_interconnect_0_data_pattern_checker_0_csr_slave_write;                       // mm_interconnect_0:data_pattern_checker_0_csr_slave_write -> data_pattern_checker_0:csr_slave_write
	wire   [31:0] mm_interconnect_0_data_pattern_checker_0_csr_slave_writedata;                   // mm_interconnect_0:data_pattern_checker_0_csr_slave_writedata -> data_pattern_checker_0:csr_slave_writedata
	wire          rst_controller_reset_out_reset;                                                 // rst_controller:reset_out -> [data_pattern_checker_0:reset_reset, data_pattern_generator_0:reset_reset, freq_counter_0:reset_n, mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset]
	wire          clk_50_clk_reset_reset;                                                         // clk_50:reset_n_out -> rst_controller:reset_in0

	xcvr_test_system_clk_50 clk_50 (
		.in_clk      (clk_50_clk),             //   input,  width = 1,       clk_in.clk
		.reset_n     (reset_50_reset_n),       //   input,  width = 1, clk_in_reset.reset_n
		.clk_out     (clk_50_clk_clk),         //  output,  width = 1,          clk.clk
		.reset_n_out (clk_50_clk_reset_reset)  //  output,  width = 1,    clk_reset.reset_n
	);

	xcvr_test_system_data_pattern_checker_0 data_pattern_checker_0 (
		.csr_clk_clk                   (clk_50_clk_clk),                                                                 //   input,    width = 1,                csr_clk.clk
		.reset_reset                   (rst_controller_reset_out_reset),                                                 //   input,    width = 1,                  reset.reset
		.csr_slave_address             (mm_interconnect_0_data_pattern_checker_0_csr_slave_address),                     //   input,    width = 3,              csr_slave.address
		.csr_slave_write               (mm_interconnect_0_data_pattern_checker_0_csr_slave_write),                       //   input,    width = 1,                       .write
		.csr_slave_read                (mm_interconnect_0_data_pattern_checker_0_csr_slave_read),                        //   input,    width = 1,                       .read
		.csr_slave_byteenable          (mm_interconnect_0_data_pattern_checker_0_csr_slave_byteenable),                  //   input,    width = 4,                       .byteenable
		.csr_slave_writedata           (mm_interconnect_0_data_pattern_checker_0_csr_slave_writedata),                   //   input,   width = 32,                       .writedata
		.csr_slave_readdata            (mm_interconnect_0_data_pattern_checker_0_csr_slave_readdata),                    //  output,   width = 32,                       .readdata
		.conduit_pattern_in_clk_export (xcvr_tx_rx_clkout2_converter_0_rx_clkout2_a_export),                             //   input,    width = 1, conduit_pattern_in_clk.export
		.asi_data                      (xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_fifo_read_export)  //   input,  width = 128,     conduit_pattern_in.export
	);

	xcvr_test_system_data_pattern_generator_0 data_pattern_generator_0 (
		.csr_clk_clk                    (clk_50_clk_clk),                                                  //   input,    width = 1,                 csr_clk.clk
		.reset_reset                    (rst_controller_reset_out_reset),                                  //   input,    width = 1,                   reset.reset
		.csr_slave_address              (mm_interconnect_0_data_pattern_generator_0_csr_slave_address),    //   input,    width = 3,               csr_slave.address
		.csr_slave_write                (mm_interconnect_0_data_pattern_generator_0_csr_slave_write),      //   input,    width = 1,                        .write
		.csr_slave_read                 (mm_interconnect_0_data_pattern_generator_0_csr_slave_read),       //   input,    width = 1,                        .read
		.csr_slave_byteenable           (mm_interconnect_0_data_pattern_generator_0_csr_slave_byteenable), //   input,    width = 4,                        .byteenable
		.csr_slave_writedata            (mm_interconnect_0_data_pattern_generator_0_csr_slave_writedata),  //   input,   width = 32,                        .writedata
		.csr_slave_readdata             (mm_interconnect_0_data_pattern_generator_0_csr_slave_readdata),   //  output,   width = 32,                        .readdata
		.conduit_pattern_out_clk_export (xcvr_tx_rx_clkout2_converter_0_tx_clkout2_a_export),              //   input,    width = 1, conduit_pattern_out_clk.export
		.aso_data                       (data_pattern_generator_0_conduit_pattern_out_export)              //  output,  width = 128,     conduit_pattern_out.export
	);

	xcvr_test_system_freq_counter_0 freq_counter_0 (
		.reset_n      (~rst_controller_reset_out_reset),                      //   input,   width = 1,        reset.reset_n
		.clk          (clk_50_clk_clk),                                       //   input,   width = 1,        clock.clk
		.csr_address  (mm_interconnect_0_freq_counter_0_csr_address),         //   input,   width = 4,          csr.address
		.csr_read     (mm_interconnect_0_freq_counter_0_csr_read),            //   input,   width = 1,             .read
		.csr_readdata (mm_interconnect_0_freq_counter_0_csr_readdata),        //  output,  width = 32,             .readdata
		.sample_clk   (xcvr_tx_rx_clkout2_converter_0_tx_clkout2_sample_clk)  //   input,   width = 1, sample_clock.clk
	);

	xcvr_test_system_mm_bridge_0 mm_bridge_0 (
		.clk              (clk_50_clk_clk),                 //   input,   width = 1,   clk.clk
		.reset            (rst_controller_reset_out_reset), //   input,   width = 1, reset.reset
		.s0_waitrequest   (mm_bridge_0_s0_waitrequest),     //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (mm_bridge_0_s0_readdata),        //  output,  width = 32,      .readdata
		.s0_readdatavalid (mm_bridge_0_s0_readdatavalid),   //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (mm_bridge_0_s0_burstcount),      //   input,   width = 1,      .burstcount
		.s0_writedata     (mm_bridge_0_s0_writedata),       //   input,  width = 32,      .writedata
		.s0_address       (mm_bridge_0_s0_address),         //   input,  width = 13,      .address
		.s0_write         (mm_bridge_0_s0_write),           //   input,   width = 1,      .write
		.s0_read          (mm_bridge_0_s0_read),            //   input,   width = 1,      .read
		.s0_byteenable    (mm_bridge_0_s0_byteenable),      //   input,   width = 4,      .byteenable
		.s0_debugaccess   (mm_bridge_0_s0_debugaccess),     //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),        //   input,  width = 32,      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),      //  output,   width = 1,      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),       //  output,  width = 32,      .writedata
		.m0_address       (mm_bridge_0_m0_address),         //  output,  width = 13,      .address
		.m0_write         (mm_bridge_0_m0_write),           //  output,   width = 1,      .write
		.m0_read          (mm_bridge_0_m0_read),            //  output,   width = 1,      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),      //  output,   width = 4,      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess)      //  output,   width = 1,      .debugaccess
	);

	xcvr_test_system_rx_fifo rx_fifo (
		.data    (xcvr_user_rx_fifo_converter_0_fifo_input_datain), //   input,   width = 64,  fifo_input.datain
		.wrreq   (xcvr_user_rx_fifo_converter_0_fifo_input_wrreq),  //   input,    width = 1,            .wrreq
		.rdreq   (xcvr_user_rx_fifo_converter_0_fifo_input_rdreq),  //   input,    width = 1,            .rdreq
		.wrclk   (xcvr_user_rx_fifo_converter_0_fifo_input_wrclk),  //   input,    width = 1,            .wrclk
		.rdclk   (xcvr_user_rx_fifo_converter_0_fifo_input_rdclk),  //   input,    width = 1,            .rdclk
		.q       (rx_fifo_fifo_output_dataout),                     //  output,  width = 128, fifo_output.dataout
		.rdempty (rx_fifo_fifo_output_rdempty),                     //  output,    width = 1,            .rdempty
		.wrfull  (rx_fifo_fifo_output_wrfull)                       //  output,    width = 1,            .wrfull
	);

	xcvr_test_system_tx_fifo tx_fifo (
		.data    (xcvr_user_tx_fifo_converter_0_fifo_input_datain), //   input,  width = 128,  fifo_input.datain
		.wrreq   (xcvr_user_tx_fifo_converter_0_fifo_input_wrreq),  //   input,    width = 1,            .wrreq
		.rdreq   (xcvr_user_tx_fifo_converter_0_fifo_input_rdreq),  //   input,    width = 1,            .rdreq
		.wrclk   (xcvr_user_tx_fifo_converter_0_fifo_input_wrclk),  //   input,    width = 1,            .wrclk
		.rdclk   (xcvr_user_tx_fifo_converter_0_fifo_input_rdclk),  //   input,    width = 1,            .rdclk
		.q       (tx_fifo_fifo_output_dataout),                     //  output,   width = 64, fifo_output.dataout
		.rdempty (tx_fifo_fifo_output_rdempty),                     //  output,    width = 1,            .rdempty
		.wrfull  (tx_fifo_fifo_output_wrfull)                       //  output,    width = 1,            .wrfull
	);

	xcvr_test_system_xcvr_tx_rx_clkout2_converter_0 xcvr_tx_rx_clkout2_converter_0 (
		.rx_clkout2        (xcvr_tx_rx_clkout2_converter_0_rx_clkout2_clk),        //   input,  width = 1,        rx_clkout2.clk
		.rx_clkout2_a      (xcvr_tx_rx_clkout2_converter_0_rx_clkout2_a_export),   //  output,  width = 1,      rx_clkout2_a.export
		.rx_clkout2_b      (xcvr_tx_rx_clkout2_converter_0_rx_clkout2_b_export),   //  output,  width = 1,      rx_clkout2_b.export
		.tx_clkout2        (xcvr_tx_rx_clkout2_converter_0_tx_clkout2_clk),        //   input,  width = 1,        tx_clkout2.clk
		.tx_clkout2_a      (xcvr_tx_rx_clkout2_converter_0_tx_clkout2_a_export),   //  output,  width = 1,      tx_clkout2_a.export
		.tx_clkout2_b      (xcvr_tx_rx_clkout2_converter_0_tx_clkout2_b_export),   //  output,  width = 1,      tx_clkout2_b.export
		.tx_clkout2_sample (xcvr_tx_rx_clkout2_converter_0_tx_clkout2_sample_clk)  //  output,  width = 1, tx_clkout2_sample.clk
	);

	xcvr_test_system_xcvr_user_rx_fifo_converter_0 xcvr_user_rx_fifo_converter_0 (
		.data_pattern_checker_pattern_in               (xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_export),           //   input,   width = 64,               data_pattern_checker_pattern_in.export
		.data_pattern_checker_pattern_in_clk           (xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_clk_export),       //   input,    width = 1,           data_pattern_checker_pattern_in_clk.export
		.data_pattern_checker_pattern_in_fifo_read     (xcvr_user_rx_fifo_converter_0_data_pattern_checker_pattern_in_fifo_read_export), //  output,  width = 128,     data_pattern_checker_pattern_in_fifo_read.export
		.data_pattern_checker_pattern_in_fifo_read_clk (xcvr_tx_rx_clkout2_converter_0_rx_clkout2_b_export),                             //   input,    width = 1, data_pattern_checker_pattern_in_fifo_read_clk.export
		.data_pattern_checker_rx_fifo_rdempty          (),                                                                               //  output,    width = 1,          data_pattern_checker_rx_fifo_rdempty.export
		.data_pattern_checker_rx_fifo_wrfull           (),                                                                               //  output,    width = 1,           data_pattern_checker_rx_fifo_wrfull.export
		.data                                          (xcvr_user_rx_fifo_converter_0_fifo_input_datain),                                //  output,   width = 64,                                    fifo_input.datain
		.wrreq                                         (xcvr_user_rx_fifo_converter_0_fifo_input_wrreq),                                 //  output,    width = 1,                                              .wrreq
		.rdreq                                         (xcvr_user_rx_fifo_converter_0_fifo_input_rdreq),                                 //  output,    width = 1,                                              .rdreq
		.wrclk                                         (xcvr_user_rx_fifo_converter_0_fifo_input_wrclk),                                 //  output,    width = 1,                                              .wrclk
		.rdclk                                         (xcvr_user_rx_fifo_converter_0_fifo_input_rdclk),                                 //  output,    width = 1,                                              .rdclk
		.q                                             (rx_fifo_fifo_output_dataout),                                                    //   input,  width = 128,                                   fifo_output.dataout
		.rdempty                                       (rx_fifo_fifo_output_rdempty),                                                    //   input,    width = 1,                                              .rdempty
		.wrfull                                        (rx_fifo_fifo_output_wrfull)                                                      //   input,    width = 1,                                              .wrfull
	);

	xcvr_test_system_xcvr_user_tx_fifo_converter_0 xcvr_user_tx_fifo_converter_0 (
		.data_pattern_generator_pattern_out                (xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_export),     //  output,   width = 64,                data_pattern_generator_pattern_out.export
		.data_pattern_generator_pattern_out_clk            (xcvr_user_tx_fifo_converter_0_data_pattern_generator_pattern_out_clk_export), //   input,    width = 1,            data_pattern_generator_pattern_out_clk.export
		.data_pattern_generator_pattern_out_fifo_write_clk (xcvr_tx_rx_clkout2_converter_0_tx_clkout2_b_export),                          //   input,    width = 1, data_pattern_generator_pattern_out_fifo_write_clk.export
		.data_pattern_generator_pattern_out_fifo_write     (data_pattern_generator_0_conduit_pattern_out_export),                         //   input,  width = 128,     data_pattern_generator_pattern_out_fifo_write.export
		.data_pattern_generator_tx_fifo_rdempty            (),                                                                            //  output,    width = 1,            data_pattern_generator_tx_fifo_rdempty.export
		.data_pattern_generator_tx_fifo_wrfull             (),                                                                            //  output,    width = 1,             data_pattern_generator_tx_fifo_wrfull.export
		.data                                              (xcvr_user_tx_fifo_converter_0_fifo_input_datain),                             //  output,  width = 128,                                        fifo_input.datain
		.wrreq                                             (xcvr_user_tx_fifo_converter_0_fifo_input_wrreq),                              //  output,    width = 1,                                                  .wrreq
		.rdreq                                             (xcvr_user_tx_fifo_converter_0_fifo_input_rdreq),                              //  output,    width = 1,                                                  .rdreq
		.wrclk                                             (xcvr_user_tx_fifo_converter_0_fifo_input_wrclk),                              //  output,    width = 1,                                                  .wrclk
		.rdclk                                             (xcvr_user_tx_fifo_converter_0_fifo_input_rdclk),                              //  output,    width = 1,                                                  .rdclk
		.q                                                 (tx_fifo_fifo_output_dataout),                                                 //   input,   width = 64,                                       fifo_output.dataout
		.rdempty                                           (tx_fifo_fifo_output_rdempty),                                                 //   input,    width = 1,                                                  .rdempty
		.wrfull                                            (tx_fifo_fifo_output_wrfull)                                                   //   input,    width = 1,                                                  .wrfull
	);

	xcvr_test_system_altera_mm_interconnect_1920_zd6ql4a mm_interconnect_0 (
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                          //   input,  width = 13,                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                                      //  output,   width = 1,                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                                       //   input,   width = 1,                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                                       //   input,   width = 4,                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                             //   input,   width = 1,                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                         //  output,  width = 32,                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                                    //  output,   width = 1,                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                            //   input,   width = 1,                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                        //   input,  width = 32,                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                                      //   input,   width = 1,                                        .debugaccess
		.freq_counter_0_csr_address                    (mm_interconnect_0_freq_counter_0_csr_address),                    //  output,   width = 4,                      freq_counter_0_csr.address
		.freq_counter_0_csr_read                       (mm_interconnect_0_freq_counter_0_csr_read),                       //  output,   width = 1,                                        .read
		.freq_counter_0_csr_readdata                   (mm_interconnect_0_freq_counter_0_csr_readdata),                   //   input,  width = 32,                                        .readdata
		.data_pattern_generator_0_csr_slave_address    (mm_interconnect_0_data_pattern_generator_0_csr_slave_address),    //  output,   width = 3,      data_pattern_generator_0_csr_slave.address
		.data_pattern_generator_0_csr_slave_write      (mm_interconnect_0_data_pattern_generator_0_csr_slave_write),      //  output,   width = 1,                                        .write
		.data_pattern_generator_0_csr_slave_read       (mm_interconnect_0_data_pattern_generator_0_csr_slave_read),       //  output,   width = 1,                                        .read
		.data_pattern_generator_0_csr_slave_readdata   (mm_interconnect_0_data_pattern_generator_0_csr_slave_readdata),   //   input,  width = 32,                                        .readdata
		.data_pattern_generator_0_csr_slave_writedata  (mm_interconnect_0_data_pattern_generator_0_csr_slave_writedata),  //  output,  width = 32,                                        .writedata
		.data_pattern_generator_0_csr_slave_byteenable (mm_interconnect_0_data_pattern_generator_0_csr_slave_byteenable), //  output,   width = 4,                                        .byteenable
		.data_pattern_checker_0_csr_slave_address      (mm_interconnect_0_data_pattern_checker_0_csr_slave_address),      //  output,   width = 3,        data_pattern_checker_0_csr_slave.address
		.data_pattern_checker_0_csr_slave_write        (mm_interconnect_0_data_pattern_checker_0_csr_slave_write),        //  output,   width = 1,                                        .write
		.data_pattern_checker_0_csr_slave_read         (mm_interconnect_0_data_pattern_checker_0_csr_slave_read),         //  output,   width = 1,                                        .read
		.data_pattern_checker_0_csr_slave_readdata     (mm_interconnect_0_data_pattern_checker_0_csr_slave_readdata),     //   input,  width = 32,                                        .readdata
		.data_pattern_checker_0_csr_slave_writedata    (mm_interconnect_0_data_pattern_checker_0_csr_slave_writedata),    //  output,  width = 32,                                        .writedata
		.data_pattern_checker_0_csr_slave_byteenable   (mm_interconnect_0_data_pattern_checker_0_csr_slave_byteenable),   //  output,   width = 4,                                        .byteenable
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                  //   input,   width = 1, mm_bridge_0_reset_reset_bridge_in_reset.reset
		.clk_50_clk_clk                                (clk_50_clk_clk)                                                   //   input,   width = 1,                              clk_50_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clk_50_clk_reset_reset),        //   input,  width = 1, reset_in0.reset
		.clk            (clk_50_clk_clk),                 //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

endmodule
